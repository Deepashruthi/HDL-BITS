module top_module();
    reg [1:0]in;
    wire out;
    
    andgate uut(.in(in), .out(out));
    
    initial begin
        in = 0;
        #10 in = 1;
        #10 in = 2;
        #10 in = 3;
        #10 $finish;
    end

endmodule
